package enum_x;

typedef enum reg[2:0] {IDLE, PHASE1, PHASE2, START, SAMPLE, SHIFT, CONTINUE} STATE;

    
endpackage