library verilog;
use verilog.vl_types.all;
entity ECL_TB is
end ECL_TB;
